`include "uvm_macros.svh"
`include "my_testbench_pkg.svh"

// The top module that contains the DUT and interface.
// This module starts the test.
module top;
    import uvm_pkg::*;
    import my_testbench_pkg::*;

    // Instantiate the interface
    dut_if dut_if1();

    // Instantiate the DUT and connect it to the interface
    dut dut1(.dif(dut_if1));

    // Clock generator
    initial begin
        dut_if1.clock = 0;
        forever #5 dut_if1.clock = ~dut_if1.clock;
    end

    initial begin
        // Place the interface into the UVM configuration database
        uvm_config_db#(virtual dut_if)::set(null, "*", "dut_vif", dut_if1);
        // Start the test
        run_test("my_test");
    end
endmodule
