`ifndef INTERF
`define INTERF

interface intf(input logic clk);
    logic [7:0] input_1;
    logic [7:0] input_2;
    logic [8:0] output_3;
endinterface
`endif 